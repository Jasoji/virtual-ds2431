library verilog;
use verilog.vl_types.all;
entity VirtualDS2431_IO_tb is
end VirtualDS2431_IO_tb;
